`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    /* Does not work with gate level sim */
    /*
    for (int i = 0; i < 35; i=i+1) $dumpvars(0, user_project.mem[i]);
    for (int i = 0; i < 16; i=i+1) $dumpvars(0, user_project.products[i]);
    for (int i = 0; i < 8; i=i+1) $dumpvars(0, user_project.sum1[i]);
    for (int i = 0; i < 4; i=i+1) $dumpvars(0, user_project.sum2[i]);
    for (int i = 0; i < 2; i=i+1) $dumpvars(0, user_project.sum3[i]);
    */
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

  // Replace tt_um_example with your module name:
  tt_um_jayjaywong12 user_project (

      // Include power ports for the Gate Level test:

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
